`ifndef ADDR_WIDTH
`define ADDR_WIDTH 32
`endif
`ifndef DATA_WIDTH
`define DATA_WIDTH 32
`endif
`ifndef NUM_WORDS
`define NUM_WORDS 16192
`endif
